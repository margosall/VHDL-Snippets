
library ieee; 
use ieee.std_logic_1164.all;

package constants is
    constant WORD_SIZE : integer := 8; -- bits for word
    constant RAM_SIZE : integer := 2; -- bits for address line
end package;


package body constants is
end constants;