
library ieee; 
use ieee.std_logic_1164.all;

package constants is
    constant SIZE : integer := 4; -- bits for input
end package;


package body constants is
end constants;