library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

PACKAGE ENC IS
	PROCEDURE SEG_CTRL (SIGNAL NUMBER : IN INTEGER RANGE 0 to 9999; SIGNAL DO0,DO1,DO2,DO3 : OUT INTEGER RANGE 0 TO 9);
END ENC;

PACKAGE BODY ENC IS
PROCEDURE SEG_CTRL (SIGNAL NUMBER : IN INTEGER RANGE 0 to 9999; SIGNAL DO0,DO1,DO2,DO3 : OUT INTEGER RANGE 0 TO 9) IS
VARIABLE TEMP: INTEGER RANGE 0 TO 9999;
VARIABLE D1: INTEGER RANGE 0 TO 9;
VARIABLE D2: INTEGER RANGE 0 TO 9;
VARIABLE D3: INTEGER RANGE 0 TO 9;
VARIABLE D4: INTEGER RANGE 0 TO 9;
BEGIN
TEMP:=NUMBER;
IF(TEMP>999) THEN
    D4:=TEMP/1000;
    TEMP:=TEMP-D4*1000;
    ELSE
    D4:=0;
END IF;
IF(TEMP > 99) THEN
    D3:=TEMP/100;
    TEMP:=TEMP-D3*100;
    ELSE
    D3:=0;
END IF;
IF(TEMP > 9) THEN
    D2:=TEMP/10;
    TEMP:=TEMP-D2*10;
    ELSE
    D2:=0;
END IF;
D1:=TEMP;

DO0<=D1;
DO1<=D2;
DO2<=D3;
DO3<=D4;
END SEG_CTRL;

END ENC;